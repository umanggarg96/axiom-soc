typedef uvm_sequencer#(apb_master_txn) apb_master_sequencer;
