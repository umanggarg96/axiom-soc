package seq_pkg;

    import uvm_pkg::*;
    import axiom_apb_pkg::*;
    `include "uvm_macros.svh"

    `include "pwm_basic_seq.svh"

endpackage
