package axiom_apb_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "master/sequence_items/apb_master_txn.svh"
    `include "master/agent/apb_master_driver.svh"
    `include "master/agent/apb_master_sequencer.svh"
    `include "master/agent/apb_master_agent.svh"
    `include "master/sequences/apb_master_base_seq.svh"

endpackage

`include "master/modules/axiom_apb_interface.sv"
`include "master/modules/axiom_apb_master.sv"
