package test_pkg;

    import uvm_pkg::*;
    import env_pkg::*;
    import seq_pkg::*;
    `include "uvm_macros.svh"

    `include "test_base.svh"

endpackage
