package seq_pkg;

    import uvm_pkg::*;
    import axiom_apb_pkg::*;
    `include "uvm_macros.svh"

    `include "uart_base_seq.svh"

endpackage
