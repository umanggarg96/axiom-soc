package env_pkg;

    import uvm_pkg::*;
    import axiom_apb_pkg::*;
    `include "uvm_macros.svh"

    `include "env.svh"

endpackage
